interface intf; 
//signal list declaration
logic [7:0] a;
logic [7:0] b;
logic [2:0] opcode;
logic [7:0] result;
logic zero;
  
endinterface
